library verilog;
use verilog.vl_types.all;
entity fakequidditch_vlg_check_tst is
    port(
        clk_out         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end fakequidditch_vlg_check_tst;
