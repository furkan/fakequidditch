library verilog;
use verilog.vl_types.all;
entity fakequidditch_vlg_vec_tst is
end fakequidditch_vlg_vec_tst;
