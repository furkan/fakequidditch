library verilog;
use verilog.vl_types.all;
entity fakequidditch is
    port(
        clk             : in     vl_logic;
        clk_out         : out    vl_logic
    );
end fakequidditch;
