module square(input number, output square);



endmodule